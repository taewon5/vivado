library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
USE ieee.std_logic_unsigned.ALL;

entity dot_matrix is 
GENERIC (clk_divider: INTEGER := 18000);    --12MHz to 500Hz
port ( rst, clk :   in std_logic;
an :   out bit_vector(7 downto 0);
dot:   out bit_vector(7 downto 0));
end dot_matrix;
-------------------------------------------------------------------
--  {0x00, 0x0e, 0x01, 0x0d, 0x13, 0x13, 0x0d,}   // 0x61, a
ARCHITECTURE dot_matrix OF dot_matrix IS
       constant N: integer :=24; -- 2^^15=32768
       TYPE state IS (S0, S1, S2, S3, S4, S5, S6, S7);
       SIGNAL pr_state, nx_state: state;
       signal r_reg, r_next: unsigned(N-1 downto 0);
       signal sel: integer:=0;
       signal     E: bit;
type Config_t is array(79 downto 0,0 to 7) of bit_vector(7 downto 0);
constant rom        : Config_t  := 
((x"00",x"00",x"04",x"08",x"1f",x"08",x"04",x"00"), -- 0x00,0x00,0x04,0x08,0x1F,0x08,0x04,0x00, <-
(x"00",x"00",x"04",x"02",x"1f",x"02",x"04",x"00"),   --0x00,0x00,0x04,0x02,0x1F,0x02,0x04,0x00, ->
(x"00",x"08",x"04",x"04",x"02",x"04",x"04",x"08"), --0x00,0x08,0x04,0x04,0x02,0x04,0x04,0x08, }
(x"00",x"04",x"04",x"04",x"04",x"04",x"04",x"04"), --0x00,0x04,0x04,0x04,0x04,0x04,0x04,0x04, |
(x"00",x"02",x"04",x"04",x"08",x"04",x"04",x"02"), --0x00,0x02,0x04,0x04,0x08,0x04,0x04,0x02, {
(x"00",x"00",x"00",x"00",x"1e",x"04",x"08",x"1e"), --0x00,0x00,0x00,0x00,0x1E,0x04,0x08,0x1E, z
(x"00",x"00",x"00",x"0a",x"0a",x"04",x"04",x"08"), -- 0x00,0x00,0x00,0x0A,0x0A,0x04,0x04,0x08, y
(x"00",x"00",x"00",x"11",x"0a",x"0a",x"0a",x"11"),   --0x00,0x00,0x00,0x11,0x0A,0x04,0x0A,0x11,x
(x"00",x"00",x"00",x"00",x"15",x"15",x"15",x"0a"), --0x00,0x00,0x00,0x00,0x15,0x15,0x15,0x0A, w
(x"00",x"00",x"00",x"00",x"14",x"14",x"14",x"08"), --0x00,0x00,0x00,0x00,0x14,0x14,0x14,0x08, v
(x"00",x"00",x"00",x"00",x"0a",x"0a",x"0a",x"0e"), --0x00,0x00,0x00,0x00,0x0A,0x0A,0x0A,0x0E, u
(x"00",x"00",x"08",x"1c",x"08",x"08",x"08",x"0c"), --0x00,0x00,0x08,0x1C,0x08,0x08,0x08,0x0C, t
(x"00",x"00",x"00",x"06",x"08",x"0e",x"02",x"0c"), --0x00,0x00,0x00,0x06,0x08,0x0E,0x02,0x0C, s
(x"00",x"00",x"00",x"0a",x"0c",x"08",x"08",x"08"), --0x00,0x00,0x00,0x0A,0x0C,0x08,0x08,0x08, r
(x"00",x"00",x"00",x"0e",x"0a",x"0e",x"02",x"02"), -- 0x00,0x00,0x00,0x0E,0x0A,0x0E,0x02,0x02, q
(x"00",x"00",x"00",x"0e",x"0a",x"0e",x"08",x"08"),   --0x00,0x00,0x00,0x0E,0x0A,0x0E,0x08,0x08, p
(x"00",x"00",x"00",x"00",x"0e",x"0a",x"0a",x"0e"), --0x00,0x00,0x00,0x00,0x0E,0x0A,0x0A,0x0E, o
(x"00",x"00",x"00",x"00",x"1e",x"12",x"12",x"12"), -- 0x00,0x00,0x00,0x00,0x1E,0x12,0x12,0x12, n
(x"00",x"00",x"00",x"11",x"1b",x"15",x"15",x"11"),  --0x00,0x00,0x00,0x11,0x1B,0x15,0x15,0x11, m
(x"00",x"00",x"04",x"04",x"04",x"04",x"04",x"04"), --0x00,0x00,0x04,0x04,0x04,0x04,0x04,0x04, l
(x"00",x"00",x"08",x"08",x"0a",x"0c",x"0a",x"0a"), -- 0x00,0x00,0x08,0x08,0x0A,0x0C,0x0A,0x0A, k
(x"00",x"00",x"04",x"00",x"04",x"04",x"04",x"08"),   --0x00,0x00,0x04,0x00,0x04,0x04,0x04,0x08,j
(x"00",x"00",x"04",x"00",x"04",x"04",x"04",x"04"), --0x00,0x00,0x04,0x00,0x04,0x04,0x04,0x04, i
(x"00",x"00",x"08",x"08",x"08",x"0e",x"0a",x"0a"), -- 0x00,0x00,0x08,0x08,0x08,0x0E,0x0A,0x0A, h
(x"00",x"0e",x"0a",x"0e",x"02",x"02",x"02",x"0e"), --0x00,0x0E,0x0A,0x0E,0x02,0x02,0x02,0x0E, g
(x"00",x"06",x"04",x"0e",x"04",x"04",x"04",x"04"), --0x00,0x06,0x04,0x0E,0x04,0x04,0x04,0x04, f
(x"00",x"00",x"00",x"04",x"0a",x"0e",x"08",x"06"), -- 0x00,0x00,0x00,0x04,0x0A,0x0E,0x08,0x06, e
(x"00",x"02",x"02",x"02",x"0e",x"12",x"12",x"0e"),  --0x00,0x02,0x02,0x02,0x0E,0x12,0x12,0x0E, d
(x"00",x"00",x"00",x"04",x"0a",x"08",x"0a",x"04"), --0x00,0x00,0x00,0x04,0x0A,0x08,0x0A,0x04, c
(x"00",x"08",x"08",x"08",x"0c",x"0a",x"0a",x"0c"), --0x00,0x08,0x08,0x08,0x0C,0x0A,0x0A,0x0C, b
(x"00",x"06",x"09",x"01",x"05",x"0a",x"0a",x"05"), --0x00,0x06,0x09,0x01,0x05,0x0A,0x0A,0x05, a
(x"00",x"08",x"04",x"02",x"00",x"00",x"00",x"00"), --0x00,0x08,0x04,0x02,0x00,0x00,0x00,0x00, `
(x"00",x"00",x"00",x"00",x"00",x"00",x"1e",x"00"), --0x00,0x00,0x00,0x00,0x00,0x00,0x1E,0x00, _
(x"00",x"04",x"0a",x"11",x"00",x"00",x"00",x"00"), --0x00,0x04,0x0A,0x11,0x00,0x00,0x00,0x00, ^
(x"00",x"00",x"0c",x"04",x"04",x"04",x"04",x"0c"), --0x00,0x00,0x0C,0x04,0x04,0x04,0x04,0x0C, ]
(x"00",x"00",x"10",x"08",x"04",x"02",x"01",x"00"), --0x00,0x00,0x10,0x08,0x04,0x02,0x01,0x00, \
(x"00",x"00",x"0c",x"08",x"08",x"08",x"08",x"0c"), --0x00,0x00,0x0C,0x08,0x08,0x08,0x08,0x0C, [
(x"00",x"1f",x"01",x"02",x"04",x"08",x"10",x"1f"),--0x00,0x1F,0x01,0x02,0x04,0x08,0x10,0x1F, Z
(x"00",x"11",x"11",x"11",x"0a",x"04",x"04",x"04"), --0x00,0x11,0x11,0x11,0x0A,0x04,0x04,0x04, Y
(x"00",x"11",x"11",x"0a",x"04",x"0a",x"11",x"11"), --0x00,0x11,0x11,0x0A,0x04,0x0A,0x11,0x11, X
(x"00",x"11",x"11",x"15",x"15",x"15",x"15",x"0a"), --0x00,0x11,0x11,0x15,0x15,0x15,0x15,0x0A, W
(x"00",x"11",x"11",x"11",x"11",x"11",x"0a",x"04"), --0x00,0x11,0x11,0x11,0x11,0x11,0x0A,0x04, V
(x"00",x"11",x"11",x"11",x"11",x"11",x"11",x"0e"),  --0x00,0x11,0x11,0x11,0x11,0x11,0x11,0x0E, U
(x"00",x"1f",x"04",x"04",x"04",x"04",x"04",x"04"), --0x00,0x1F,0x04,0x04,0x04,0x04,0x04,0x04, T
(x"00",x"0e",x"10",x"10",x"1e",x"02",x"02",x"1c"), --0x00,0x0E,0x10,0x10,0x1E,0x02,0x02,0x1C, S
(x"00",x"0c",x"12",x"12",x"1e",x"18",x"14",x"12"), --0x00,0x1C,0x12,0x12,0x1E,0x18,0x14,0x12, R
(x"00",x"0c",x"12",x"12",x"12",x"12",x"14",x"0a"), --0x00,0x0C,0x12,0x12,0x12,0x12,0x14,0x0A, Q
(x"00",x"1c",x"12",x"12",x"1c",x"10",x"10",x"10"), --0x00,0x1C,0x12,0x12,0x1C,0x10,0x10,0x10, P
(x"00",x"0e",x"11",x"11",x"11",x"11",x"11",x"0e"), --0x00,0x0E,0x11,0x11,0x11,0x11,0x11,0x0E, O
(x"00",x"11",x"11",x"19",x"15",x"13",x"11",x"11"), --0x00,0x11,0x11,0x19,0x15,0x13,0x11,0x11, N
(x"00",x"11",x"1b",x"15",x"15",x"11",x"11",x"11"), --0x00,0x11,0x1B,0x15,0x15,0x11,0x11,0x11, M
(x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"1e"), --0x00,0x10,0x10,0x10,0x10,0x10,0x10,0x1E, L 
(x"00",x"11",x"12",x"14",x"18",x"14",x"12",x"11"), --0x00,0x11,0x12,0x14,0x18,0x14,0x12,0x11, K
(x"00",x"02",x"02",x"02",x"02",x"12",x"12",x"0c"), --0x00,0x02,0x02,0x02,0x02,0x12,0x12,0x0C, J
(x"00",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c"), --0x00,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C,0x0C, I
(x"00",x"12",x"12",x"12",x"1e",x"12",x"12",x"12"), --0x00,0x12,0x12,0x12,0x1E,0x12,0x12,0x12, H
(x"00",x"0c",x"12",x"10",x"16",x"12",x"12",x"0c"), --0x00,0x0C,0x12,0x10,0x16,0x12,0x12,0x0C, G
(x"00",x"1e",x"10",x"10",x"1e",x"10",x"10",x"10"), --0x00,0x1E,0x10,0x10,0x1E,0x10,0x10,0x10, F
(x"00",x"1e",x"10",x"10",x"1e",x"10",x"10",x"1e"), -- 0x00,0x1E,0x10,0x10,0x1E,0x10,0x10,0x1E, E
(x"00",x"1c",x"12",x"12",x"12",x"12",x"1c",x"00"),  --0x00,0x1C,0x12,0x12,0x12,0x12,0x1C,0x00, D
(x"00",x"0c",x"12",x"10",x"10",x"10",x"12",x"0c"), --0x00,0x0C,0x12,0x10,0x10,0x10,0x12,0x0C,, C
(x"1c",x"12",x"12",x"1c",x"12",x"12",x"1c",x"00"), --0x1C,0x12,0x12,0x1C,0x12,0x12,0x1C,0x00, B
(x"0e",x"0e",x"11",x"11",x"1f",x"11",x"11",x"11"), --0x00,0x0E,0x11,0x11,0x1F,0x11,0x11,0x11, A
(x"0e",x"11",x"01",x"0d",x"15",x"15",x"0e",x"00"), --0x0E,0x11,0x01,0x0D,0x15,0x15,0x0E,0x00, @
(x"0e",x"11",x"01",x"02",x"04",x"00",x"04",x"00"), --0x0E,0x11,0x01,0x02,0x04,0x00,0x04,0x00, ?
(x"00",x"10",x"08",x"04",x"02",x"04",x"08",x"10"), --0x00,0x10,0x08,0x04,0x02,0x04,0x08,0x10,>
(x"00",x"00",x"1e",x"00",x"1e",x"00",x"00",x"00"), --0x00,0x00,0x1E,0x00,0x1E,0x00,0x00,0x00, =
(x"00",x"02",x"04",x"08",x"10",x"08",x"04",x"02"), --0x00,0x02,0x04,0x08,0x10,0x08,0x04,0x02, <
(x"00",x"0c",x"0c",x"00",x"00",x"0c",x"04",x"08"), --0x00,0x0C,0x0C,0x00,0x00,0x0C,0x04,0x08, ;
(x"00",x"0c",x"0c",x"00",x"00",x"0c",x"0c",x"00"), --0x00,0x0C,0x0C,0x00,0x00,0x0C,0x0C,0x00, :
(x"00",x"0c",x"12",x"12",x"0e",x"02",x"12",x"0c"), --0x00,0x0C,0x12,0x12,0x0E,0x02,0x12,0x0C, 9
(x"00",x"1e",x"12",x"12",x"1e",x"12",x"12",x"1e"), --0x00,0x1E,0x12,0x12,0x1E,0x12,0x12,0x1E, 8
(x"00",x"1e",x"12",x"12",x"02",x"02",x"02",x"02"), --0x00,0x1E,0x12,0x12,0x02,0x02,0x02,0x02, 7
(x"00",x"0c",x"12",x"10",x"1c",x"12",x"12",x"0c"), --0x00,0x0C,0x12,0x10,0x1C,0x12,0x12,0x0C, 6
(x"00",x"1e",x"10",x"10",x"0c",x"02",x"02",x"1c"), --0x00,0x1E,0x10,0x10,0x0C,0x02,0x02,0x1C, 5
(x"02",x"06",x"0a",x"12",x"1f",x"02",x"02",x"00"), --0x02,0x06,0x0A,0x12,0x1F,0x02,0x02,0x00,4
(x"00",x"0c",x"12",x"02",x"0e",x"02",x"12",x"0c"), --0x00,0x0C,0x12,0x02,0x0E,0x02,0x12,0x0C, 3
(x"0c",x"1e",x"12",x"02",x"04",x"08",x"10",x"1e"),--0x0C,0x1E,0x12,0x02,0x04,0x08,0x10,0x1E, 2
(x"04",x"0c",x"1c",x"0c",x"0c",x"0c",x"0c",x"1e"), --0x04,0x0C,0x1C,0x0C,0x0C,0x0C,0x0C,0x1E, 1
(x"00",x"0c",x"12",x"12",x"16",x"1a",x"12",x"0c") --0x00,0x0C,0x12,0x12,0x16,0x1A,0x12,0x0C, 0 
                                        );
BEGIN
----- Clock generator (E->500Hz): -------------
PROCESS (clk)
VARIABLE count: INTEGER RANGE 0 TO clk_divider;
BEGIN
IF (clk'EVENT AND clk='1') THEN
count := count + 1;
IF (count=clk_divider) THEN
E <= NOT E;
count := 0;
 END IF;
END IF;
END PROCESS;
 ----- Lower section of FSM: --------------------
PROCESS (E)
BEGIN
 IF (E'EVENT AND E='1') THEN
 IF (rst='1') THEN
  pr_state <= S0;
ELSE
 pr_state <= nx_state;
 END IF;
 END IF;
 END PROCESS;
 
process(clk)
begin
if(clk'event and clk='1') then
r_reg <= r_next;
if(r_reg="111111111111111111111111") then
sel<=sel + 1;
end if;
end if;
end process;
r_next <= r_reg + 1;


PROCESS (sel,pr_state)
 BEGIN
-- register
 CASE pr_state IS
  WHEN S0 =>
  dot<=rom(sel,0);
  an <= "01111111";
  nx_state <= S1;
 WHEN S1 =>
  dot<=rom(sel,1);
  an <= "10111111";
  nx_state <= S2;
 WHEN S2 =>
  dot<=rom(sel,2);
  an <= "11011111";
  nx_state <= S3;
   WHEN S3 =>
    dot<=rom(sel,3);
   an <= "11101111";
     nx_state <= S4;
    WHEN S4 =>
  dot<=rom(sel,4);
  an <= "11110111";
  nx_state <= S5;
   WHEN S5 =>
   dot<=rom(sel,5);
  an <= "11111011";
    nx_state <= S6;
  WHEN S6 =>
     dot<=rom(sel,6);
      an <= "11111101";
       nx_state <= S7;
    WHEN S7 =>
       dot<=rom(sel,7);
       an <= "11111110";
       nx_state <= S0;
   END CASE;
   END PROCESS;
END dot_matrix;